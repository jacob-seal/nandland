-- Package file containing all Constants and Components used in Pong Game

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package Pong_Pkg is

  -----------------------------------------------------------------------------
  -- Constants
  -----------------------------------------------------------------------------
  
  -- Set the Width and Height of the Game Board
  constant c_Game_Width    : integer := 40;
  constant c_Game_Height   : integer := 30;

  -- Set the number of points to play to
  constant c_Score_Limit : integer := 5;
  
  -- Set the Height (in board game units) of the paddle.
  constant c_Paddle_Height : integer := 6;

  -- Set the Speed of the paddle movement.  In this case, the paddle will move
  -- one board game unit every 50 milliseconds that the button is held down.
  constant c_Paddle_Speed : integer := 1250000;

  -- Set the Speed of the ball movement.  In this case, the ball will move
  -- one board game unit every 50 milliseconds that the button is held down.   
  constant c_Ball_Speed : integer  := 2500000;
  
  -- Sets Column index to draw Player 1 & Player 2 Paddles.
  constant c_Paddle_Col_Location_P1 : integer := 0;
  constant c_Paddle_Col_Location_P2 : integer := c_Game_Width-1;

  --constants for score offset
  constant c_x_offset_p1 : integer := 230;
  constant c_x_offset_p2 : integer := 390;
  constant c_y_offset_p1_p2 : integer := 10;

  -----------------------------------------------------------------------------
  -- Numeric bit patterns for output to VGA for scorekeeping
  -----------------------------------------------------------------------------
  type bitmap_type is array (0 to 19) of std_logic_vector(0 to 49);
	-- '0'
  constant c_zero_bmp : bitmap_type := 
    (
        ("00000000000000000000000000000000000000000000000000"),
        ("00000000000000000000000000000000000000000000000000"),
        ("00000000000001111111111111111111111100000000000000"),
        ("00000000000001110000000000000000011100000000000000"),
        ("00000000000001110000000000000000011100000000000000"),
        ("00000000000001110000000000000000011100000000000000"),
        ("00000000000001110000000000000000011100000000000000"),
        ("00000000000001110000000000000000011100000000000000"),
        ("00000000000001110000000000000000011100000000000000"),
        ("00000000000001110000000000000000011100000000000000"),
        ("00000000000001110000000000000000011100000000000000"),
        ("00000000000001110000000000000000011100000000000000"),
        ("00000000000001110000000000000000011100000000000000"),
        ("00000000000001110000000000000000011100000000000000"),
        ("00000000000001110000000000000000011100000000000000"),
        ("00000000000001110000000000000000011100000000000000"),
        ("00000000000001110000000000000000011100000000000000"),
        ("00000000000001111111111111111111111100000000000000"),
        ("00000000000000000000000000000000000000000000000000"),
        ("00000000000000000000000000000000000000000000000000")
    );
  -- '1'
  constant c_one_bmp : bitmap_type := 
    (
        ("00000000000000000000000000000000000000000000000000"),
        ("00000000000000000000000000000000000000000000000000"),
        ("00000000000000000000111111000000000000000000000000"),
        ("00000000000000000011111111000000000000000000000000"),
        ("00000000000000000000000111000000000000000000000000"),
        ("00000000000000000000000111000000000000000000000000"),
        ("00000000000000000000000111000000000000000000000000"),
        ("00000000000000000000000111000000000000000000000000"),
        ("00000000000000000000000111000000000000000000000000"),
        ("00000000000000000000000111000000000000000000000000"),
        ("00000000000000000000000111000000000000000000000000"),
        ("00000000000000000000000111000000000000000000000000"),
        ("00000000000000000000000111000000000000000000000000"),
        ("00000000000000000000000111000000000000000000000000"),
        ("00000000000000000000000111000000000000000000000000"),
        ("00000000000000000000000111000000000000000000000000"),
        ("00000000000000000111111111111111000000000000000000"),
        ("00000000000000000111111111111111000000000000000000"),
        ("00000000000000000000000000000000000000000000000000"),
        ("00000000000000000000000000000000000000000000000000")
    );
    -- '2'
  constant c_two_bmp : bitmap_type := 
    (
        ("00000000000000000000000000000000000000000000000000"),
        ("00000000000000000000000000000000000000000000000000"),
        ("00000000000001111111111111111111100000000000000000"),
        ("00000000000001111111111111111111100000000000000000"),
        ("00000000000000000000000000000011100000000000000000"),
        ("00000000000000000000000000000011100000000000000000"),
        ("00000000000000000000000000000011100000000000000000"),
        ("00000000000000000000000000000011100000000000000000"),
        ("00000000000000000000000000000011100000000000000000"),
        ("00000000000001111111111111111111100000000000000000"),
        ("00000000000001111111111111111111100000000000000000"),
        ("00000000000001110000000000000000000000000000000000"),
        ("00000000000001110000000000000000000000000000000000"),
        ("00000000000001110000000000000000000000000000000000"),
        ("00000000000001110000000000000000000000000000000000"),
        ("00000000000001110000000000000000000000000000000000"),
        ("00000000000001111111111111111111100000000000000000"),
        ("00000000000001111111111111111111100000000000000000"),
        ("00000000000000000000000000000000000000000000000000"),
        ("00000000000000000000000000000000000000000000000000")
    );
    -- '3'
  constant c_three_bmp : bitmap_type := 
    (
        ("00000000000000000000000000000000000000000000000000"),
        ("00000000000000000000000000000000000000000000000000"),
        ("00000000000001111111111111111111100000000000000000"),
        ("00000000000001111111111111111111100000000000000000"),
        ("00000000000000000000000000000011100000000000000000"),
        ("00000000000000000000000000000011100000000000000000"),
        ("00000000000000000000000000000011100000000000000000"),
        ("00000000000000000000000000000011100000000000000000"),
        ("00000000000000000000000000000011100000000000000000"),
        ("00000000000000000111111111111111100000000000000000"),
        ("00000000000000000111111111111111100000000000000000"),
        ("00000000000000000000000000000011100000000000000000"),
        ("00000000000000000000000000000011100000000000000000"),
        ("00000000000000000000000000000011100000000000000000"),
        ("00000000000000000000000000000011100000000000000000"),
        ("00000000000000000000000000000011100000000000000000"),
        ("00000000000001111111111111111111100000000000000000"),
        ("00000000000001111111111111111111100000000000000000"),
        ("00000000000000000000000000000000000000000000000000"),
        ("00000000000000000000000000000000000000000000000000")
    );
    -- '4'
  constant c_four_bmp : bitmap_type := 
    (
        ("00000000000000000000000000000000000000000000000000"),
        ("00000000000000000000000000000000000000000000000000"),
        ("00000000000001110000000000000000111000000000000000"),
        ("00000000000001110000000000000000111000000000000000"),
        ("00000000000001110000000000000000111000000000000000"),
        ("00000000000001110000000000000000111000000000000000"),
        ("00000000000001110000000000000000111000000000000000"),
        ("00000000000001110000000000000000111000000000000000"),
        ("00000000000001110000000000000000111000000000000000"),
        ("00000000000001111111111111111111111000000000000000"),
        ("00000000000001111111111111111111111000000000000000"),
        ("00000000000000000000000000000000111000000000000000"),
        ("00000000000000000000000000000000111000000000000000"),
        ("00000000000000000000000000000000111000000000000000"),
        ("00000000000000000000000000000000111000000000000000"),
        ("00000000000000000000000000000000111000000000000000"),
        ("00000000000000000000000000000000111000000000000000"),
        ("00000000000000000000000000000000111000000000000000"),
        ("00000000000000000000000000000000000000000000000000"),
        ("00000000000000000000000000000000000000000000000000")
    );
    -- '5'
  constant c_five_bmp : bitmap_type := 
    (
        ("00000000000000000000000000000000000000000000000000"),
        ("00000000000000000000000000000000000000000000000000"),
        ("00000000000001111111111111111111111000000000000000"),
        ("00000000000001111111111111111111111000000000000000"),
        ("00000000000001110000000000000000000000000000000000"),
        ("00000000000001110000000000000000000000000000000000"),
        ("00000000000001110000000000000000000000000000000000"),
        ("00000000000001110000000000000000000000000000000000"),
        ("00000000000001110000000000000000000000000000000000"),
        ("00000000000001111111111111111111111000000000000000"),
        ("00000000000001111111111111111111111000000000000000"),
        ("00000000000000000000000000000000111000000000000000"),
        ("00000000000000000000000000000000111000000000000000"),
        ("00000000000000000000000000000000111000000000000000"),
        ("00000000000000000000000000000000111000000000000000"),
        ("00000000000000000000000000000000111000000000000000"),
        ("00000000000001111111111111111111111000000000000000"),
        ("00000000000001111111111111111111111000000000000000"),
        ("00000000000000000000000000000000000000000000000000"),
        ("00000000000000000000000000000000000000000000000000")
    );


  -----------------------------------------------------------------------------
  -- Component Declarations
  -----------------------------------------------------------------------------
  component Pong_Paddle_Ctrl is
    generic (
      g_Player_Paddle_X : integer  -- Changes for P1 vs P2
      );
    port (
      i_Clk : in std_logic;

      i_Col_Count_Div : in std_logic_vector(5 downto 0);
      i_Row_Count_Div : in std_logic_vector(5 downto 0);

      -- Player Paddle Control
      i_Paddle_Up : in std_logic;
      i_Paddle_Dn : in std_logic;

      o_Draw_Paddle : out std_logic;
      o_Paddle_Y    : out std_logic_vector(5 downto 0)
      );
  end component Pong_Paddle_Ctrl;


  component Pong_Ball_Ctrl is
    port (
      i_Clk           : in  std_logic;
      i_Game_Active   : in  std_logic;
      i_Col_Count_Div : in  std_logic_vector(5 downto 0);
      i_Row_Count_Div : in  std_logic_vector(5 downto 0);
      --
      o_Draw_Ball     : out std_logic;
      o_Ball_X        : out std_logic_vector(5 downto 0);
      o_Ball_Y        : out std_logic_vector(5 downto 0)
      );
  end component Pong_Ball_Ctrl;

  
  component Pong_Score_Ctrl is
    generic (
    g_X_offset : integer  -- Changes for P1 vs P2
    );
    port (
      i_Clk           : in std_logic;
      i_score         : in integer;
      i_Col_Count     : in std_logic_vector(9 downto 0);
      i_Row_Count     : in std_logic_vector(9 downto 0);
      o_Draw_Score   : out std_logic
      );
  end component Pong_Score_Ctrl;  


  
end package Pong_Pkg;  
